module alu(

);